// -*- Verilog -*-


`define DIFFTEST
//  `define SIMUTEST
// `define BTB_LOG
// `define BTB_CLOSE
`define BIG_CACHE
`define UNCACHE
// `define IBAR
//`define OURDIV