module EX2_WB(
    
);
endmodule