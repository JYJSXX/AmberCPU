// -*- Verilog -*-

`ifdef VERILATOR
`define CONFIG_DIFFTEST
// `define CONFIG_BR_PROFILE
// `define CONFIG_INST_PROFILE
// `define CONFIG_AXI_PROFILE
// `define CONFIG_LD_ST_PROFILE
// `define CONFIG_CACHE_PROFILE
`endif
