
module TLB(
    
);

endmodule