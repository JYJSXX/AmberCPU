module IQ (
    // TODO Dispatch
);
    
endmodule