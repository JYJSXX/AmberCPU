module moduleName (
    input [31:0]        inst0_i,
    input [31:0]        inst1_i,
    output [3:0]        type_
);
    
endmodule