module EX_Privilege(
    input clk,
    input rstn,

    input en,
    input csr,
    input [31:0] rd_data,
    input [31:0] rj_data,
    input [13:0] csr_num,
    
);

endmodule