// `include "define.vh"
// module BTB_local (
//     input           clk,
//     input           rstn,
//     input   [31:0]  fact_tpc,
//     input           fact_taken,
//     output          pred_taken
// );
//     wire [7:0] HASH_INDEX;
//     reg  [];

//     assign      HASH_INDEX  =   {fact_tpc[17:13],fact_tpc[5:3]};

// endmodule