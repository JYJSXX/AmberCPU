`include "../config.vh"
`include "../exception.vh"

module TLB_EXP(
    input [31:0] vaddr0,
    input en0,
    input [1:0] plv0, //crmd_plv
    input is_if_0,
    input is_store_0,
    input is_load_0,
    

    input [31:0] vaddr1,
);
endmodule