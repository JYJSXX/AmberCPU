// -*- Verilog -*-


`define DIFFTEST
// `define SIMUTEST
// `define BTB_LOG
`define BTB_CLOSE
// `define BR_PROFILE
// `define INST_PROFILE
// `define AXI_PROFILE
// `define LD_ST_PROFILE
// `define CACHE_PROFILE

